module RBLut(
		output[15:0] lut[4:0]
	);
	
	assign lut = '{16'd23};
endmodule
