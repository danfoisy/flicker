// FrameBuf_single.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module FrameBuf_single (
		input  wire        clk_clk,       //   clk.clk
		input  wire        reset_reset,   // reset.reset
		input  wire [11:0] s1_address,    //    s1.address
		input  wire        s1_clken,      //      .clken
		input  wire        s1_chipselect, //      .chipselect
		input  wire        s1_write,      //      .write
		output wire [15:0] s1_readdata,   //      .readdata
		input  wire [15:0] s1_writedata,  //      .writedata
		input  wire [1:0]  s1_byteenable  //      .byteenable
	);

	FrameBuf_single_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),       //   clk1.clk
		.address    (s1_address),    //     s1.address
		.clken      (s1_clken),      //       .clken
		.chipselect (s1_chipselect), //       .chipselect
		.write      (s1_write),      //       .write
		.readdata   (s1_readdata),   //       .readdata
		.writedata  (s1_writedata),  //       .writedata
		.byteenable (s1_byteenable), //       .byteenable
		.reset      (reset_reset),   // reset1.reset
		.reset_req  (1'b0),          // (terminated)
		.freeze     (1'b0)           // (terminated)
	);

endmodule
