// FrameBuf_lg.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module FrameBuf_lg (
		input  wire        mem_clk1_clk,      // mem_clk1.clk
		input  wire        mem_clk2_clk,      // mem_clk2.clk
		input  wire        mem_rst1_reset,    // mem_rst1.reset
		input  wire        mem_rst2_reset,    // mem_rst2.reset
		input  wire [13:0] mem_s1_address,    //   mem_s1.address
		input  wire        mem_s1_clken,      //         .clken
		input  wire        mem_s1_chipselect, //         .chipselect
		input  wire        mem_s1_write,      //         .write
		output wire [15:0] mem_s1_readdata,   //         .readdata
		input  wire [15:0] mem_s1_writedata,  //         .writedata
		input  wire [1:0]  mem_s1_byteenable, //         .byteenable
		input  wire [13:0] mem_s2_address,    //   mem_s2.address
		input  wire        mem_s2_chipselect, //         .chipselect
		input  wire        mem_s2_clken,      //         .clken
		input  wire        mem_s2_write,      //         .write
		output wire [15:0] mem_s2_readdata,   //         .readdata
		input  wire [15:0] mem_s2_writedata,  //         .writedata
		input  wire [1:0]  mem_s2_byteenable  //         .byteenable
	);

	FrameBuf_lg_onchip_memory2_0 onchip_memory2_0 (
		.clk         (mem_clk1_clk),      //   clk1.clk
		.address     (mem_s1_address),    //     s1.address
		.clken       (mem_s1_clken),      //       .clken
		.chipselect  (mem_s1_chipselect), //       .chipselect
		.write       (mem_s1_write),      //       .write
		.readdata    (mem_s1_readdata),   //       .readdata
		.writedata   (mem_s1_writedata),  //       .writedata
		.byteenable  (mem_s1_byteenable), //       .byteenable
		.reset       (mem_rst1_reset),    // reset1.reset
		.address2    (mem_s2_address),    //     s2.address
		.chipselect2 (mem_s2_chipselect), //       .chipselect
		.clken2      (mem_s2_clken),      //       .clken
		.write2      (mem_s2_write),      //       .write
		.readdata2   (mem_s2_readdata),   //       .readdata
		.writedata2  (mem_s2_writedata),  //       .writedata
		.byteenable2 (mem_s2_byteenable), //       .byteenable
		.clk2        (mem_clk2_clk),      //   clk2.clk
		.reset2      (mem_rst2_reset),    // reset2.reset
		.reset_req   (1'b0),              // (terminated)
		.freeze      (1'b0),              // (terminated)
		.reset_req2  (1'b0)               // (terminated)
	);

endmodule
